// (c) Technion IIT, Department of Electrical Engineering 2018 

// Implements a simple equality one-bit out comparator
// with a parameter Nbits to define the inputs' size


module comparator 
	(
   // Input, Output Ports
	input logic [3:0] vect1,
	input logic [3:0] vect2,
	output logic cmp
   );
	
   assign cmp = (vect1 == vect2);

endmodule
