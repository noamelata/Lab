
module	gameoverBMP (
					 
					output	logic	[0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors  //rgb value from the bitmap 
 ) ;
 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 6;  // 2^6 = 64 
localparam  int OBJECT_NUMBER_OF_X_BITS = 6;  // 2^6 = 64 


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

assign object_colors = {
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff, 8'hff, 8'hff, 8'hff, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff },
{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff }
};


endmodule