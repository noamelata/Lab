

module GAME_TOP	(	
					input		logic	clk,
					input		logic	resetN,
					
					input		logic	playerDrawingRequest,	
					input		logic	[7:0] treesDrawingRequest,			
					output	logic SingleHitPulse
					
);
endmodule

