
module	heartBMP (
					 
					output	logic	[0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_color  //rgb value from the bitmap 
 ) ;
 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^5 = 32 


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

assign object_color = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hFA, 8'hFA, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hFF, 8'hFF, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hFF, 8'hFF },
{8'hFF, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hFA, 8'hFA, 8'hFA, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hFF },
{8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hE9, 8'hE9, 8'hE9, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hE9, 8'hE9, 8'hE9, 8'hFA, 8'hFA, 8'hFA, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hC9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hC9, 8'hC9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hC9, 8'hC9, 8'hC9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4 },
{8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF },
{8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hA4, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA4, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};


endmodule